`timescale 1ns/1ps  //时间精度
`define    Clock 20 //时钟周期

module FSM_3_tb;
//--------------------< 端口 >------------------------------------------
reg                     clk                 ;
reg                     rst_n               ;
reg  [1:0]              in                  ;
wire [1:0]              out                 ;
wire                    out_vld             ;

//----------------------------------------------------------------------
//--   模块例化
//----------------------------------------------------------------------
FSM_3 u_FSM_3
(
    .clk                (clk                ),
    .rst_n              (rst_n              ),
    .in                 (in                 ),
    .out                (out                ),
    .out_vld            (out_vld            )
);

//----------------------------------------------------------------------
//--   状态机名称查看器
//----------------------------------------------------------------------
localparam S0           = 4'b0001           ;
localparam S1           = 4'b0010           ;
localparam S2           = 4'b0100           ;
localparam S3           = 4'b1000           ;
//2字符16位
reg [15:0]              state_name          ;

always@(*)begin
    case(u_FSM_3.state_c)
        S0:     state_name = "S0";
        S1:     state_name = "S1";
        S2:     state_name = "S2";
        S3:     state_name = "S3";
        default:state_name = "S0";
    endcase
end

//----------------------------------------------------------------------
//--   时钟信号和复位信号
//----------------------------------------------------------------------
initial begin
    clk = 1;
    forever
    #(`Clock/2) clk = ~clk;
end

initial begin
    rst_n = 0; #(`Clock*20+1);
    rst_n = 1;
end

//----------------------------------------------------------------------
//--   设计输入信号
//----------------------------------------------------------------------
initial begin

    $dumpfile("test.vcd");
    $dumpvars(0,FSM_3_tb);
    #1;
    in = 0;
    #(`Clock*20+1); //初始化完成
//情况1--------------------------
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*10);
//情况2--------------------------
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*10);
//情况3--------------------------
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*10);
//情况4--------------------------
    in = 1;         //1块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*10);
//情况5--------------------------
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*1);
    in = 2;         //2块钱
    #(`Clock*1);
    in = 0;
    #(`Clock*10);


    $stop;
end


endmodule

